// +FHDR--------------------------------------------------------------------------------------------
// Copyright (c) 2016 Xxx.
// -------------------------------------------------------------------------------------------------
// Filename      : alu.v
// Author        : r04099
// Created On    : 2016-01-11 23:47
// Last Modified : 2016-01-11 23:47
// -------------------------------------------------------------------------------------------------
// Svn Info:
//   $Revision::                                                                                $:
//   $Author::                                                                                  $:
//   $Date::                                                                                    $:
//   $HeadURL::                                                                                 $:
// -------------------------------------------------------------------------------------------------
// Description:
//
//
// -FHDR--------------------------------------------------------------------------------------------

module alu ( a, b, cmd, r );
  input [15:0] a;
  input [15:0] b;
  input [2:0] cmd;
  output [15:0] r;
  wire   \C4/DATA8_0 , \C4/DATA8_1 , \C4/DATA8_2 , \C4/DATA8_3 , \C4/DATA8_4 ,
         \C4/DATA8_5 , \C4/DATA8_6 , \C4/DATA8_7 , \C4/DATA8_8 , \C4/DATA8_9 ,
         \C4/DATA8_10 , \C4/DATA8_11 , \C4/DATA8_12 , \C4/DATA8_13 ,
         \C4/DATA8_14 , \DP_OP_21J1_124_1250/n53 , \DP_OP_21J1_124_1250/n36 ,
         \DP_OP_21J1_124_1250/n35 , \DP_OP_21J1_124_1250/n34 ,
         \DP_OP_21J1_124_1250/n33 , \DP_OP_21J1_124_1250/n32 ,
         \DP_OP_21J1_124_1250/n31 , \DP_OP_21J1_124_1250/n30 ,
         \DP_OP_21J1_124_1250/n29 , \DP_OP_21J1_124_1250/n28 ,
         \DP_OP_21J1_124_1250/n27 , \DP_OP_21J1_124_1250/n26 ,
         \DP_OP_21J1_124_1250/n25 , \DP_OP_21J1_124_1250/n24 ,
         \DP_OP_21J1_124_1250/n23 , \DP_OP_21J1_124_1250/n22 ,
         \DP_OP_21J1_124_1250/n16 , \DP_OP_21J1_124_1250/n15 ,
         \DP_OP_21J1_124_1250/n14 , \DP_OP_21J1_124_1250/n13 ,
         \DP_OP_21J1_124_1250/n12 , \DP_OP_21J1_124_1250/n11 ,
         \DP_OP_21J1_124_1250/n10 , \DP_OP_21J1_124_1250/n9 ,
         \DP_OP_21J1_124_1250/n8 , \DP_OP_21J1_124_1250/n7 ,
         \DP_OP_21J1_124_1250/n6 , \DP_OP_21J1_124_1250/n5 ,
         \DP_OP_21J1_124_1250/n4 , \DP_OP_21J1_124_1250/n3 ,
         \DP_OP_21J1_124_1250/n2 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347;

  ADDFXL \DP_OP_21J1_124_1250/U17  ( .A(a[0]), .B(\DP_OP_21J1_124_1250/n53 ), 
        .CI(\DP_OP_21J1_124_1250/n36 ), .CO(\DP_OP_21J1_124_1250/n16 ), .S(
        \C4/DATA8_0 ) );
  ADDFXL \DP_OP_21J1_124_1250/U16  ( .A(\DP_OP_21J1_124_1250/n35 ), .B(a[1]), 
        .CI(\DP_OP_21J1_124_1250/n16 ), .CO(\DP_OP_21J1_124_1250/n15 ), .S(
        \C4/DATA8_1 ) );
  ADDFXL \DP_OP_21J1_124_1250/U15  ( .A(\DP_OP_21J1_124_1250/n34 ), .B(a[2]), 
        .CI(\DP_OP_21J1_124_1250/n15 ), .CO(\DP_OP_21J1_124_1250/n14 ), .S(
        \C4/DATA8_2 ) );
  ADDFXL \DP_OP_21J1_124_1250/U14  ( .A(\DP_OP_21J1_124_1250/n33 ), .B(a[3]), 
        .CI(\DP_OP_21J1_124_1250/n14 ), .CO(\DP_OP_21J1_124_1250/n13 ), .S(
        \C4/DATA8_3 ) );
  ADDFXL \DP_OP_21J1_124_1250/U13  ( .A(\DP_OP_21J1_124_1250/n32 ), .B(a[4]), 
        .CI(\DP_OP_21J1_124_1250/n13 ), .CO(\DP_OP_21J1_124_1250/n12 ), .S(
        \C4/DATA8_4 ) );
  ADDFXL \DP_OP_21J1_124_1250/U12  ( .A(\DP_OP_21J1_124_1250/n31 ), .B(a[5]), 
        .CI(\DP_OP_21J1_124_1250/n12 ), .CO(\DP_OP_21J1_124_1250/n11 ), .S(
        \C4/DATA8_5 ) );
  ADDFXL \DP_OP_21J1_124_1250/U10  ( .A(\DP_OP_21J1_124_1250/n29 ), .B(a[7]), 
        .CI(\DP_OP_21J1_124_1250/n10 ), .CO(\DP_OP_21J1_124_1250/n9 ), .S(
        \C4/DATA8_7 ) );
  ADDFXL \DP_OP_21J1_124_1250/U8  ( .A(\DP_OP_21J1_124_1250/n27 ), .B(a[9]), 
        .CI(\DP_OP_21J1_124_1250/n8 ), .CO(\DP_OP_21J1_124_1250/n7 ), .S(
        \C4/DATA8_9 ) );
  ADDFXL \DP_OP_21J1_124_1250/U7  ( .A(\DP_OP_21J1_124_1250/n26 ), .B(a[10]), 
        .CI(\DP_OP_21J1_124_1250/n7 ), .CO(\DP_OP_21J1_124_1250/n6 ), .S(
        \C4/DATA8_10 ) );
  ADDFXL \DP_OP_21J1_124_1250/U6  ( .A(\DP_OP_21J1_124_1250/n25 ), .B(a[11]), 
        .CI(\DP_OP_21J1_124_1250/n6 ), .CO(\DP_OP_21J1_124_1250/n5 ), .S(
        \C4/DATA8_11 ) );
  ADDFXL \DP_OP_21J1_124_1250/U5  ( .A(\DP_OP_21J1_124_1250/n24 ), .B(a[12]), 
        .CI(\DP_OP_21J1_124_1250/n5 ), .CO(\DP_OP_21J1_124_1250/n4 ), .S(
        \C4/DATA8_12 ) );
  ADDFXL \DP_OP_21J1_124_1250/U4  ( .A(\DP_OP_21J1_124_1250/n23 ), .B(a[13]), 
        .CI(\DP_OP_21J1_124_1250/n4 ), .CO(\DP_OP_21J1_124_1250/n3 ), .S(
        \C4/DATA8_13 ) );
  XOR2XL \DP_OP_21J1_124_1250/U35  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[0]), 
        .Y(\DP_OP_21J1_124_1250/n36 ) );
  XOR2XL \DP_OP_21J1_124_1250/U34  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[1]), 
        .Y(\DP_OP_21J1_124_1250/n35 ) );
  XOR2XL \DP_OP_21J1_124_1250/U30  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[5]), 
        .Y(\DP_OP_21J1_124_1250/n31 ) );
  XOR2XL \DP_OP_21J1_124_1250/U31  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[4]), 
        .Y(\DP_OP_21J1_124_1250/n32 ) );
  XOR2XL \DP_OP_21J1_124_1250/U32  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[3]), 
        .Y(\DP_OP_21J1_124_1250/n33 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U33  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[2]), 
        .Y(\DP_OP_21J1_124_1250/n34 ) );
  ADDFXL \DP_OP_21J1_124_1250/U9  ( .A(\DP_OP_21J1_124_1250/n28 ), .B(a[8]), 
        .CI(\DP_OP_21J1_124_1250/n9 ), .CO(\DP_OP_21J1_124_1250/n8 ), .S(
        \C4/DATA8_8 ) );
  ADDFXL \DP_OP_21J1_124_1250/U3  ( .A(\DP_OP_21J1_124_1250/n22 ), .B(a[14]), 
        .CI(\DP_OP_21J1_124_1250/n3 ), .CO(\DP_OP_21J1_124_1250/n2 ), .S(
        \C4/DATA8_14 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U27  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[8]), 
        .Y(\DP_OP_21J1_124_1250/n28 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U28  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[7]), 
        .Y(\DP_OP_21J1_124_1250/n29 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U29  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[6]), 
        .Y(\DP_OP_21J1_124_1250/n30 ) );
  ADDFXL \DP_OP_21J1_124_1250/U11  ( .A(\DP_OP_21J1_124_1250/n30 ), .B(a[6]), 
        .CI(\DP_OP_21J1_124_1250/n11 ), .CO(\DP_OP_21J1_124_1250/n10 ), .S(
        \C4/DATA8_6 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U26  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[9]), 
        .Y(\DP_OP_21J1_124_1250/n27 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U25  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[10]), 
        .Y(\DP_OP_21J1_124_1250/n26 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U24  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[11]), 
        .Y(\DP_OP_21J1_124_1250/n25 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U23  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[12]), 
        .Y(\DP_OP_21J1_124_1250/n24 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U22  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[13]), 
        .Y(\DP_OP_21J1_124_1250/n23 ) );
  XOR2X1 \DP_OP_21J1_124_1250/U21  ( .A(\DP_OP_21J1_124_1250/n53 ), .B(b[14]), 
        .Y(\DP_OP_21J1_124_1250/n22 ) );
  OAI22XL U2 ( .A0(b[1]), .A1(n160), .B0(n190), .B1(n292), .Y(n1) );
  OAI21XL U3 ( .A0(n42), .A1(n1), .B0(n180), .Y(n338) );
  NOR2BX1 U4 ( .AN(n69), .B(n72), .Y(\DP_OP_21J1_124_1250/n53 ) );
  AOI222XL U5 ( .A0(n210), .A1(n129), .B0(b[1]), .B1(n189), .C0(n211), .C1(
        n310), .Y(n2) );
  OAI22XL U6 ( .A0(n284), .A1(n308), .B0(n326), .B1(n2), .Y(n3) );
  OAI21XL U7 ( .A0(n324), .A1(n238), .B0(n273), .Y(n4) );
  OAI22XL U8 ( .A0(b[0]), .A1(n41), .B0(n343), .B1(n272), .Y(n5) );
  OAI211X1 U9 ( .A0(n329), .A1(n309), .B0(n331), .C0(n5), .Y(n6) );
  CLKINVX1 U10 ( .A(n308), .Y(n7) );
  NAND2X1 U11 ( .A(n211), .B(a[0]), .Y(n8) );
  OAI211X1 U12 ( .A0(n190), .A1(n189), .B0(n83), .C0(n8), .Y(n9) );
  AO22X1 U13 ( .A0(b[2]), .A1(n238), .B0(n42), .B1(n9), .Y(n10) );
  NOR2X1 U14 ( .A(n305), .B(n10), .Y(n11) );
  AOI211X1 U15 ( .A0(n176), .A1(n7), .B0(n287), .C0(n11), .Y(n12) );
  OAI21XL U16 ( .A0(n332), .A1(a[0]), .B0(n331), .Y(n13) );
  AO22X1 U17 ( .A0(b[0]), .A1(n13), .B0(n69), .B1(\C4/DATA8_0 ), .Y(n14) );
  AOI211X1 U18 ( .A0(a[0]), .A1(n6), .B0(n12), .C0(n14), .Y(n15) );
  OAI31XL U19 ( .A0(n262), .A1(n3), .A2(n4), .B0(n15), .Y(r[0]) );
  OAI21XL U20 ( .A0(n284), .A1(n274), .B0(n273), .Y(n16) );
  OAI21XL U21 ( .A0(n326), .A1(n276), .B0(n298), .Y(n17) );
  AOI211X1 U22 ( .A0(n275), .A1(n277), .B0(n16), .C0(n17), .Y(n18) );
  OAI2BB2XL U23 ( .B0(n42), .B1(n277), .A0N(n42), .A1N(n276), .Y(n19) );
  OAI2BB2XL U24 ( .B0(n305), .B1(n19), .A0N(n278), .A1N(n279), .Y(n20) );
  AOI211X1 U25 ( .A0(b[3]), .A1(n280), .B0(n287), .C0(n20), .Y(n21) );
  AOI211X1 U26 ( .A0(n281), .A1(n313), .B0(n18), .C0(n21), .Y(n22) );
  OAI21XL U27 ( .A0(n332), .A1(b[6]), .B0(n331), .Y(n23) );
  AOI22X1 U28 ( .A0(a[6]), .A1(n23), .B0(n69), .B1(\C4/DATA8_6 ), .Y(n24) );
  AO22X1 U29 ( .A0(a[6]), .A1(n272), .B0(n271), .B1(n41), .Y(n25) );
  OAI21XL U30 ( .A0(n317), .A1(n25), .B0(b[6]), .Y(n26) );
  NAND3X1 U31 ( .A(n22), .B(n24), .C(n26), .Y(r[6]) );
  OAI22XL U32 ( .A0(n309), .A1(n346), .B0(n332), .B1(b[15]), .Y(n27) );
  AOI211X1 U33 ( .A0(n272), .A1(b[15]), .B0(n317), .C0(n27), .Y(n28) );
  AOI2BB2X1 U34 ( .B0(\DP_OP_21J1_124_1250/n53 ), .B1(b[15]), .A0N(
        \DP_OP_21J1_124_1250/n53 ), .A1N(b[15]), .Y(n29) );
  AOI2BB2X1 U35 ( .B0(a[15]), .B1(n29), .A0N(a[15]), .A1N(n29), .Y(n30) );
  AOI2BB2X1 U36 ( .B0(\DP_OP_21J1_124_1250/n2 ), .B1(n30), .A0N(
        \DP_OP_21J1_124_1250/n2 ), .A1N(n30), .Y(n31) );
  OAI21XL U37 ( .A0(a[15]), .A1(n332), .B0(n331), .Y(n32) );
  AO22X1 U38 ( .A0(n69), .A1(n31), .B0(b[15]), .B1(n32), .Y(n33) );
  AOI31X1 U39 ( .A0(n253), .A1(n155), .A2(n285), .B0(n33), .Y(n34) );
  CLKINVX1 U40 ( .A(n156), .Y(n35) );
  OAI21XL U41 ( .A0(n330), .A1(n303), .B0(n329), .Y(n36) );
  OAI22XL U42 ( .A0(a[14]), .A1(n215), .B0(a[15]), .B1(n170), .Y(n37) );
  OAI22XL U43 ( .A0(n213), .A1(a[13]), .B0(n214), .B1(a[12]), .Y(n38) );
  OAI21XL U44 ( .A0(n37), .A1(n38), .B0(n296), .Y(n39) );
  OAI211X1 U45 ( .A0(n324), .A1(n35), .B0(n36), .C0(n39), .Y(n40) );
  OAI211X1 U46 ( .A0(n292), .A1(n28), .B0(n34), .C0(n40), .Y(r[15]) );
  CLKINVX1 U47 ( .A(b[2]), .Y(n42) );
  OAI31XL U48 ( .A0(n287), .A1(n206), .A2(n205), .B0(n204), .Y(r[2]) );
  AOI211X1 U49 ( .A0(n306), .A1(n274), .B0(n151), .C0(n150), .Y(n152) );
  AOI211X1 U50 ( .A0(n191), .A1(a[8]), .B0(n89), .C0(n88), .Y(n147) );
  AOI211X1 U51 ( .A0(n339), .A1(n338), .B0(n337), .C0(n336), .Y(n341) );
  AOI211X1 U52 ( .A0(a[6]), .A1(n193), .B0(n166), .C0(n164), .Y(n125) );
  OAI211X1 U53 ( .A0(n300), .A1(n299), .B0(n298), .C0(n297), .Y(n301) );
  NOR3X1 U54 ( .A(n293), .B(n292), .C(n309), .Y(n299) );
  AOI211X1 U55 ( .A0(n295), .A1(n288), .B0(n287), .C0(n286), .Y(n290) );
  NAND2X1 U56 ( .A(b[2]), .B(n339), .Y(n283) );
  AOI211X1 U57 ( .A0(n258), .A1(n339), .B0(n287), .C0(n257), .Y(n260) );
  NOR3X1 U58 ( .A(b[2]), .B(n193), .C(n292), .Y(n254) );
  NAND2X1 U59 ( .A(n190), .B(n42), .Y(n124) );
  OAI211X1 U60 ( .A0(n247), .A1(n305), .B0(n246), .C0(n245), .Y(n248) );
  OAI211X1 U61 ( .A0(n241), .A1(n284), .B0(n240), .C0(n340), .Y(n242) );
  AOI211X1 U62 ( .A0(n275), .A1(n239), .B0(n262), .C0(n233), .Y(n236) );
  NOR2X1 U63 ( .A(n293), .B(n231), .Y(n232) );
  AOI32XL U64 ( .A0(a[15]), .A1(b[2]), .A2(n211), .B0(n294), .B1(n42), .Y(n225) );
  AOI211X1 U65 ( .A0(\C4/DATA8_3 ), .A1(n69), .B0(n56), .C0(n55), .Y(n229) );
  AOI211X1 U66 ( .A0(n279), .A1(n220), .B0(n287), .C0(n219), .Y(n223) );
  OAI211X1 U67 ( .A0(a[5]), .A1(n213), .B0(n42), .C0(n212), .Y(n217) );
  NAND2X1 U68 ( .A(n273), .B(n82), .Y(n330) );
  AOI211X1 U69 ( .A0(\C4/DATA8_1 ), .A1(n69), .B0(n52), .C0(n51), .Y(n185) );
  AOI211X1 U70 ( .A0(n191), .A1(n221), .B0(b[2]), .C0(n171), .Y(n172) );
  NOR2XL U71 ( .A(b[4]), .B(b[3]), .Y(n339) );
  NAND2X1 U72 ( .A(n300), .B(n82), .Y(n329) );
  NOR2XL U73 ( .A(cmd[1]), .B(n78), .Y(n82) );
  NOR2XL U74 ( .A(b[3]), .B(n293), .Y(n300) );
  NAND2XL U75 ( .A(n70), .B(cmd[1]), .Y(n321) );
  NOR2X1 U76 ( .A(cmd[2]), .B(cmd[1]), .Y(n69) );
  NOR2XL U77 ( .A(n42), .B(b[3]), .Y(n275) );
  NOR2XL U78 ( .A(b[3]), .B(b[2]), .Y(n296) );
  INVXL U79 ( .A(cmd[0]), .Y(n72) );
  INVXL U80 ( .A(cmd[2]), .Y(n70) );
  INVXL U81 ( .A(cmd[1]), .Y(n71) );
  NOR2XL U82 ( .A(b[4]), .B(n81), .Y(n273) );
  NOR4XL U83 ( .A(b[13]), .B(b[8]), .C(n77), .D(n76), .Y(n246) );
  INVXL U84 ( .A(b[3]), .Y(n284) );
  NOR2X1 U85 ( .A(n214), .B(n292), .Y(n75) );
  INVXL U86 ( .A(a[15]), .Y(n292) );
  NOR2XL U87 ( .A(n190), .B(b[0]), .Y(n191) );
  NOR2XL U88 ( .A(n343), .B(b[1]), .Y(n210) );
  INVXL U89 ( .A(b[0]), .Y(n343) );
  INVXL U90 ( .A(b[1]), .Y(n190) );
  AOI211X1 U91 ( .A0(\C4/DATA8_2 ), .A1(n69), .B0(n54), .C0(n53), .Y(n204) );
  AND2X2 U92 ( .A(a[2]), .B(n196), .Y(n54) );
  OAI211X1 U93 ( .A0(n153), .A1(n154), .B0(n152), .C0(n67), .Y(n68) );
  NAND2X1 U94 ( .A(a[14]), .B(n137), .Y(n67) );
  AOI211X1 U95 ( .A0(n288), .A1(n278), .B0(n149), .C0(n280), .Y(n150) );
  OAI211X1 U96 ( .A0(a[12]), .A1(n213), .B0(n145), .C0(n144), .Y(n146) );
  NAND2X1 U97 ( .A(n211), .B(n143), .Y(n144) );
  NAND2X1 U98 ( .A(n141), .B(n281), .Y(n148) );
  CLKINVX1 U99 ( .A(a[14]), .Y(n143) );
  CLKINVX1 U100 ( .A(b[14]), .Y(n153) );
  AOI211X1 U101 ( .A0(\C4/DATA8_13 ), .A1(n69), .B0(n50), .C0(n49), .Y(n136)
         );
  OAI211X1 U102 ( .A0(n324), .A1(n325), .B0(n131), .C0(n130), .Y(n132) );
  AND2X2 U103 ( .A(b[13]), .B(n135), .Y(n50) );
  OAI211X1 U104 ( .A0(n346), .A1(n231), .B0(n122), .C0(n121), .Y(r[12]) );
  OAI211X1 U105 ( .A0(n311), .A1(n324), .B0(n120), .C0(n119), .Y(n121) );
  AOI211X1 U106 ( .A0(\C4/DATA8_12 ), .A1(n69), .B0(n48), .C0(n47), .Y(n122)
         );
  AOI211X1 U107 ( .A0(n244), .A1(n288), .B0(n109), .C0(n149), .Y(n111) );
  CLKINVX1 U108 ( .A(n307), .Y(n149) );
  AND2X2 U109 ( .A(b[12]), .B(n112), .Y(n48) );
  OAI211X1 U110 ( .A0(n346), .A1(n225), .B0(n108), .C0(n107), .Y(r[11]) );
  OAI211X1 U111 ( .A0(n294), .A1(n195), .B0(n307), .C0(n218), .Y(n107) );
  CLKINVX1 U112 ( .A(n288), .Y(n195) );
  AOI211X1 U113 ( .A0(\C4/DATA8_11 ), .A1(n69), .B0(n46), .C0(n45), .Y(n108)
         );
  NOR4X1 U114 ( .A(n102), .B(n101), .C(n165), .D(n167), .Y(n156) );
  NOR2X1 U115 ( .A(n213), .B(n322), .Y(n101) );
  AND2X2 U116 ( .A(b[11]), .B(n106), .Y(n46) );
  OAI211X1 U117 ( .A0(n199), .A1(n346), .B0(n96), .C0(n95), .Y(r[10]) );
  OAI211X1 U118 ( .A0(n305), .A1(n194), .B0(n307), .C0(n342), .Y(n95) );
  AOI211X1 U119 ( .A0(\C4/DATA8_10 ), .A1(n69), .B0(n44), .C0(n43), .Y(n96) );
  NAND2X1 U120 ( .A(n141), .B(n200), .Y(n90) );
  NOR2X1 U121 ( .A(b[2]), .B(n139), .Y(n200) );
  CLKINVX1 U122 ( .A(n330), .Y(n141) );
  AND2X2 U123 ( .A(b[10]), .B(n93), .Y(n44) );
  OAI211X1 U124 ( .A0(n347), .A1(n346), .B0(n345), .C0(n344), .Y(r[9]) );
  OAI211X1 U125 ( .A0(n343), .A1(n342), .B0(n341), .C0(n340), .Y(n344) );
  CLKINVX1 U126 ( .A(n155), .Y(n337) );
  AOI211X1 U127 ( .A0(\C4/DATA8_9 ), .A1(n69), .B0(n64), .C0(n63), .Y(n345) );
  AND2X2 U128 ( .A(b[9]), .B(n335), .Y(n64) );
  CLKINVX1 U129 ( .A(n306), .Y(n346) );
  OAI211X1 U130 ( .A0(n303), .A1(n329), .B0(n302), .C0(n301), .Y(r[7]) );
  AOI211X1 U131 ( .A0(\C4/DATA8_7 ), .A1(n69), .B0(n62), .C0(n61), .Y(n302) );
  NOR2X1 U132 ( .A(n305), .B(b[2]), .Y(n288) );
  AND2X2 U133 ( .A(b[7]), .B(n291), .Y(n62) );
  AOI211X1 U134 ( .A0(a[5]), .A1(n191), .B0(n209), .C0(n100), .Y(n157) );
  AOI211X1 U135 ( .A0(a[9]), .A1(n193), .B0(n187), .C0(n186), .Y(n188) );
  NOR2X1 U136 ( .A(n213), .B(n315), .Y(n186) );
  NOR2X1 U137 ( .A(b[2]), .B(n138), .Y(n274) );
  AOI211X1 U138 ( .A0(a[12]), .A1(n191), .B0(n80), .C0(n79), .Y(n277) );
  NOR2X1 U139 ( .A(n170), .B(n207), .Y(n80) );
  AOI21X1 U140 ( .A0(n211), .A1(a[2]), .B0(n84), .Y(n139) );
  AOI211X1 U141 ( .A0(a[4]), .A1(n191), .B0(n187), .C0(n86), .Y(n140) );
  NOR2X1 U142 ( .A(n170), .B(n271), .Y(n187) );
  OAI211X1 U143 ( .A0(n270), .A1(n329), .B0(n269), .C0(n268), .Y(r[5]) );
  OAI211X1 U144 ( .A0(n267), .A1(n326), .B0(n266), .C0(n265), .Y(n268) );
  NAND2X1 U145 ( .A(n275), .B(n264), .Y(n265) );
  NAND2X1 U146 ( .A(n42), .B(n181), .Y(n263) );
  AOI211X1 U147 ( .A0(\C4/DATA8_5 ), .A1(n69), .B0(n60), .C0(n59), .Y(n269) );
  CLKINVX1 U148 ( .A(n252), .Y(n267) );
  AND2X2 U149 ( .A(b[5]), .B(n261), .Y(n60) );
  OAI211X1 U150 ( .A0(n221), .A1(n213), .B0(n128), .C0(n169), .Y(n323) );
  CLKINVX1 U151 ( .A(a[4]), .Y(n192) );
  OAI211X1 U152 ( .A0(n250), .A1(n329), .B0(n249), .C0(n248), .Y(r[4]) );
  AOI211X1 U153 ( .A0(n244), .A1(n279), .B0(n243), .C0(n242), .Y(n245) );
  AOI211X1 U154 ( .A0(\C4/DATA8_4 ), .A1(n69), .B0(n58), .C0(n57), .Y(n249) );
  NAND2BX1 U155 ( .AN(n244), .B(n42), .Y(n231) );
  AND2X2 U156 ( .A(a[4]), .B(n235), .Y(n58) );
  AOI32X1 U157 ( .A0(a[0]), .A1(b[2]), .A2(n211), .B0(n42), .B1(n314), .Y(n250) );
  OAI211X1 U158 ( .A0(n230), .A1(n329), .B0(n229), .C0(n228), .Y(r[3]) );
  CLKINVX1 U159 ( .A(n220), .Y(n294) );
  NAND2X1 U160 ( .A(n211), .B(n221), .Y(n212) );
  AOI211X1 U161 ( .A0(a[8]), .A1(n210), .B0(n209), .C0(n208), .Y(n295) );
  NOR2X1 U162 ( .A(n170), .B(n282), .Y(n209) );
  CLKINVX1 U163 ( .A(n241), .Y(n109) );
  NOR2X1 U164 ( .A(n102), .B(n97), .Y(n220) );
  NOR2X1 U165 ( .A(n170), .B(n162), .Y(n102) );
  NOR2X1 U166 ( .A(b[2]), .B(n255), .Y(n279) );
  NOR2X1 U167 ( .A(n222), .B(n284), .Y(n56) );
  NAND2X1 U168 ( .A(n42), .B(n158), .Y(n230) );
  OAI211X1 U169 ( .A0(n129), .A1(n213), .B0(n99), .C0(n98), .Y(n158) );
  NAND2X1 U170 ( .A(n193), .B(a[0]), .Y(n98) );
  NAND4X1 U171 ( .A(n319), .B(n318), .C(n320), .D(n65), .Y(n66) );
  NAND2X1 U172 ( .A(a[8]), .B(n304), .Y(n65) );
  NOR2X1 U173 ( .A(n287), .B(n336), .Y(n307) );
  OAI211X1 U174 ( .A0(n215), .A1(n282), .B0(n114), .C0(n113), .Y(n311) );
  CLKINVX1 U175 ( .A(a[5]), .Y(n251) );
  NOR3X1 U176 ( .A(n310), .B(n309), .C(n330), .Y(n312) );
  CLKINVX1 U177 ( .A(n329), .Y(n313) );
  OAI211X1 U178 ( .A0(n129), .A1(n214), .B0(n116), .C0(n115), .Y(n314) );
  OAI211X1 U179 ( .A0(n328), .A1(n329), .B0(n185), .C0(n184), .Y(r[1]) );
  AOI211X1 U180 ( .A0(n176), .A1(n338), .B0(n287), .C0(n175), .Y(n178) );
  NAND2X1 U181 ( .A(b[2]), .B(n193), .Y(n174) );
  CLKINVX1 U182 ( .A(a[3]), .Y(n221) );
  NOR4BX1 U183 ( .AN(n169), .B(n168), .C(n167), .D(n166), .Y(n252) );
  NOR2X1 U184 ( .A(n213), .B(n282), .Y(n166) );
  CLKINVX1 U185 ( .A(a[7]), .Y(n282) );
  NOR2X1 U186 ( .A(n214), .B(n315), .Y(n167) );
  CLKINVX1 U187 ( .A(a[8]), .Y(n315) );
  NOR2X1 U188 ( .A(n215), .B(n271), .Y(n168) );
  CLKINVX1 U189 ( .A(a[6]), .Y(n271) );
  NAND2X1 U190 ( .A(n211), .B(a[5]), .Y(n169) );
  NAND2X1 U191 ( .A(n264), .B(n42), .Y(n180) );
  NOR3X1 U192 ( .A(n165), .B(n164), .C(n163), .Y(n264) );
  NOR2X1 U193 ( .A(n170), .B(n322), .Y(n164) );
  NOR2X1 U194 ( .A(n215), .B(n207), .Y(n165) );
  AND2X2 U195 ( .A(a[1]), .B(n177), .Y(n52) );
  NAND2X1 U196 ( .A(n159), .B(n42), .Y(n328) );
  NAND2X1 U197 ( .A(n155), .B(n340), .Y(n287) );
  NOR2X1 U198 ( .A(n81), .B(n243), .Y(n155) );
  CLKINVX1 U199 ( .A(n339), .Y(n305) );
  NAND2X1 U200 ( .A(n210), .B(a[1]), .Y(n83) );
  CLKINVX1 U201 ( .A(n255), .Y(n176) );
  CLKINVX1 U202 ( .A(n321), .Y(n272) );
  CLKINVX1 U203 ( .A(n332), .Y(n41) );
  NAND2X1 U204 ( .A(n211), .B(n42), .Y(n309) );
  CLKINVX1 U205 ( .A(n273), .Y(n293) );
  CLKINVX1 U206 ( .A(n317), .Y(n331) );
  NOR2X1 U207 ( .A(n72), .B(n321), .Y(n317) );
  NAND3X1 U208 ( .A(n71), .B(n72), .C(cmd[2]), .Y(n332) );
  NAND4X1 U209 ( .A(n115), .B(n113), .C(n85), .D(n87), .Y(n238) );
  NAND2X1 U210 ( .A(n193), .B(a[7]), .Y(n87) );
  NAND2X1 U211 ( .A(n210), .B(a[5]), .Y(n85) );
  NAND2X1 U212 ( .A(n191), .B(a[6]), .Y(n113) );
  NAND2X1 U213 ( .A(n211), .B(a[4]), .Y(n115) );
  CLKINVX1 U214 ( .A(n275), .Y(n324) );
  CLKINVX1 U215 ( .A(n296), .Y(n326) );
  CLKINVX1 U216 ( .A(a[0]), .Y(n310) );
  CLKINVX1 U217 ( .A(a[1]), .Y(n129) );
  CLKINVX1 U218 ( .A(n298), .Y(n262) );
  NOR3X1 U219 ( .A(n71), .B(n70), .C(n72), .Y(n298) );
  NAND2X1 U220 ( .A(n246), .B(n240), .Y(n81) );
  CLKINVX1 U221 ( .A(b[5]), .Y(n240) );
  AOI211X1 U222 ( .A0(a[14]), .A1(n191), .B0(n75), .C0(n74), .Y(n244) );
  CLKINVX1 U223 ( .A(a[12]), .Y(n161) );
  CLKINVX1 U224 ( .A(a[13]), .Y(n142) );
  AOI211X1 U225 ( .A0(n211), .A1(a[8]), .B0(n89), .C0(n73), .Y(n239) );
  CLKINVX1 U226 ( .A(a[11]), .Y(n162) );
  CLKINVX1 U227 ( .A(n193), .Y(n214) );
  NOR2X1 U228 ( .A(n190), .B(n343), .Y(n193) );
  CLKINVX1 U229 ( .A(a[10]), .Y(n207) );
  CLKINVX1 U230 ( .A(n191), .Y(n213) );
  NOR2X1 U231 ( .A(n215), .B(n322), .Y(n89) );
  CLKINVX1 U232 ( .A(a[9]), .Y(n322) );
  CLKINVX1 U233 ( .A(n210), .Y(n215) );
  CLKINVX1 U234 ( .A(n170), .Y(n211) );
  NAND2X1 U235 ( .A(n190), .B(n343), .Y(n170) );
  AO21X1 U236 ( .A0(b[2]), .A1(n203), .B0(n202), .Y(n53) );
  AOI211XL U237 ( .A0(n199), .A1(b[3]), .B0(n293), .C0(n198), .Y(n201) );
  AO21X1 U238 ( .A0(n69), .A1(\C4/DATA8_14 ), .B0(n68), .Y(r[14]) );
  AO21X1 U239 ( .A0(a[13]), .A1(n123), .B0(n134), .Y(n49) );
  AO21X1 U240 ( .A0(a[12]), .A1(n110), .B0(n111), .Y(n47) );
  AO21X1 U241 ( .A0(a[11]), .A1(n104), .B0(n105), .Y(n45) );
  AO21X1 U242 ( .A0(a[10]), .A1(n91), .B0(n92), .Y(n43) );
  NAND3XL U243 ( .A(b[4]), .B(b[2]), .C(b[1]), .Y(n342) );
  AO21X1 U244 ( .A0(a[9]), .A1(n333), .B0(n334), .Y(n63) );
  AO21X1 U245 ( .A0(a[7]), .A1(n289), .B0(n290), .Y(n61) );
  AOI21XL U246 ( .A0(b[4]), .A1(n309), .B0(n292), .Y(n285) );
  AOI211XL U247 ( .A0(b[3]), .A1(n263), .B0(n293), .C0(n262), .Y(n266) );
  AO21X1 U248 ( .A0(a[5]), .A1(n259), .B0(n260), .Y(n59) );
  AO21X1 U249 ( .A0(b[4]), .A1(n237), .B0(n236), .Y(n57) );
  AOI211XL U250 ( .A0(b[3]), .A1(n225), .B0(n293), .C0(n262), .Y(n226) );
  AO21X1 U251 ( .A0(a[3]), .A1(n224), .B0(n223), .Y(n55) );
  AO21X1 U252 ( .A0(n69), .A1(\C4/DATA8_8 ), .B0(n66), .Y(r[8]) );
  AOI211XL U253 ( .A0(b[3]), .A1(n347), .B0(n293), .C0(n262), .Y(n182) );
  AO21X1 U254 ( .A0(b[1]), .A1(n179), .B0(n178), .Y(n51) );
  NAND2XL U255 ( .A(b[4]), .B(b[3]), .Y(n253) );
  NAND2XL U256 ( .A(b[4]), .B(n292), .Y(n340) );
  NAND3XL U257 ( .A(cmd[2]), .B(cmd[1]), .C(n72), .Y(n243) );
  NAND2XL U258 ( .A(n234), .B(b[3]), .Y(n255) );
  INVXL U259 ( .A(b[4]), .Y(n234) );
  NAND2XL U260 ( .A(cmd[2]), .B(cmd[0]), .Y(n78) );
  OAI22XL U261 ( .A0(n213), .A1(n207), .B0(n214), .B1(n162), .Y(n73) );
  OAI22XL U262 ( .A0(n215), .A1(n142), .B0(n170), .B1(n161), .Y(n74) );
  OAI22XL U263 ( .A0(b[2]), .A1(n239), .B0(n42), .B1(n244), .Y(n308) );
  OR4X1 U264 ( .A(b[10]), .B(b[12]), .C(b[15]), .D(b[11]), .Y(n77) );
  OR4X1 U265 ( .A(b[14]), .B(b[6]), .C(b[9]), .D(b[7]), .Y(n76) );
  OAI22XL U266 ( .A0(b[0]), .A1(a[2]), .B0(n343), .B1(a[3]), .Y(n189) );
  OAI221XL U267 ( .A0(b[0]), .A1(a[14]), .B0(n343), .B1(a[15]), .C0(n190), .Y(
        n138) );
  OAI22XL U268 ( .A0(n214), .A1(n142), .B0(n215), .B1(n162), .Y(n79) );
  OR2X1 U269 ( .A(n277), .B(b[2]), .Y(n94) );
  OA21XL U270 ( .A0(n42), .A1(n138), .B0(n94), .Y(n199) );
  NOR3X1 U271 ( .A(n262), .B(n81), .C(n305), .Y(n306) );
  OAI221XL U272 ( .A0(a[10]), .A1(n332), .B0(n207), .B1(n321), .C0(n331), .Y(
        n93) );
  OAI21XL U273 ( .A0(n310), .A1(n213), .B0(n83), .Y(n84) );
  OAI21XL U274 ( .A0(n221), .A1(n214), .B0(n85), .Y(n86) );
  OAI21XL U275 ( .A0(n207), .A1(n170), .B0(n87), .Y(n88) );
  AOI222XL U276 ( .A0(n90), .A1(n329), .B0(n275), .B1(n140), .C0(n296), .C1(
        n147), .Y(n92) );
  OAI21XL U277 ( .A0(b[10]), .A1(n332), .B0(n331), .Y(n91) );
  OAI22XL U278 ( .A0(n211), .A1(a[15]), .B0(n170), .B1(a[14]), .Y(n278) );
  OAI21XL U279 ( .A0(n42), .A1(n278), .B0(n94), .Y(n194) );
  OAI21XL U280 ( .A0(a[15]), .A1(n284), .B0(n253), .Y(n336) );
  OAI22XL U281 ( .A0(b[0]), .A1(a[13]), .B0(n343), .B1(a[14]), .Y(n160) );
  OAI22XL U282 ( .A0(n160), .A1(n190), .B0(n215), .B1(n161), .Y(n97) );
  OAI221XL U283 ( .A0(a[11]), .A1(n332), .B0(n162), .B1(n321), .C0(n331), .Y(
        n106) );
  AOI2BB2X1 U284 ( .B0(n210), .B1(a[2]), .A0N(n170), .A1N(n221), .Y(n99) );
  OR2X1 U285 ( .A(n230), .B(n330), .Y(n103) );
  OAI22XL U286 ( .A0(n214), .A1(n192), .B0(n215), .B1(n271), .Y(n100) );
  AOI222XL U287 ( .A0(n103), .A1(n329), .B0(n275), .B1(n157), .C0(n296), .C1(
        n156), .Y(n105) );
  OAI21XL U288 ( .A0(b[11]), .A1(n332), .B0(n331), .Y(n104) );
  OAI21XL U289 ( .A0(n292), .A1(b[4]), .B0(b[2]), .Y(n241) );
  OAI21XL U290 ( .A0(n170), .A1(n292), .B0(n109), .Y(n218) );
  OAI221XL U291 ( .A0(a[12]), .A1(n332), .B0(n161), .B1(n321), .C0(n331), .Y(
        n112) );
  OAI21XL U292 ( .A0(b[12]), .A1(n332), .B0(n331), .Y(n110) );
  AOI2BB2X1 U293 ( .B0(n211), .B1(a[8]), .A0N(n214), .A1N(n251), .Y(n114) );
  AOI2BB2X1 U294 ( .B0(n191), .B1(a[2]), .A0N(n215), .A1N(n221), .Y(n116) );
  OAI21XL U295 ( .A0(n250), .A1(n330), .B0(n329), .Y(n120) );
  OAI22XL U296 ( .A0(a[12]), .A1(n170), .B0(a[11]), .B1(n215), .Y(n118) );
  OAI22XL U297 ( .A0(a[10]), .A1(n213), .B0(a[9]), .B1(n214), .Y(n117) );
  OAI21XL U298 ( .A0(n118), .A1(n117), .B0(n296), .Y(n119) );
  OAI22XL U299 ( .A0(b[1]), .A1(n160), .B0(n292), .B1(n213), .Y(n181) );
  OAI221XL U300 ( .A0(a[13]), .A1(n332), .B0(n142), .B1(n321), .C0(n331), .Y(
        n135) );
  OAI21XL U301 ( .A0(b[13]), .A1(n332), .B0(n331), .Y(n123) );
  OAI2BB2XL U302 ( .B0(n160), .B1(n124), .A0N(a[15]), .A1N(n124), .Y(n256) );
  OAI22XL U303 ( .A0(n256), .A1(n305), .B0(n254), .B1(n234), .Y(n133) );
  OAI21XL U304 ( .A0(n215), .A1(n315), .B0(n125), .Y(n325) );
  OAI22XL U305 ( .A0(a[13]), .A1(n170), .B0(a[12]), .B1(n215), .Y(n127) );
  OAI22XL U306 ( .A0(a[10]), .A1(n214), .B0(a[11]), .B1(n213), .Y(n126) );
  OAI21XL U307 ( .A0(n127), .A1(n126), .B0(n296), .Y(n131) );
  AOI2BB2X1 U308 ( .B0(n193), .B1(a[2]), .A0N(n215), .A1N(n192), .Y(n128) );
  AOI221XL U309 ( .A0(b[0]), .A1(n310), .B0(n343), .B1(n129), .C0(b[1]), .Y(
        n159) );
  OAI22XL U310 ( .A0(b[2]), .A1(n323), .B0(n42), .B1(n159), .Y(n270) );
  OAI21XL U311 ( .A0(n270), .A1(n330), .B0(n329), .Y(n130) );
  OAI31XL U312 ( .A0(n336), .A1(n337), .A2(n133), .B0(n132), .Y(n134) );
  OAI21XL U313 ( .A0(n346), .A1(n263), .B0(n136), .Y(r[13]) );
  AOI221XL U314 ( .A0(n272), .A1(a[14]), .B0(n41), .B1(n143), .C0(n317), .Y(
        n154) );
  OAI21XL U315 ( .A0(b[14]), .A1(n332), .B0(n331), .Y(n137) );
  OAI22XL U316 ( .A0(b[2]), .A1(n140), .B0(n42), .B1(n139), .Y(n281) );
  AOI2BB2X1 U317 ( .B0(n210), .B1(n142), .A0N(n214), .A1N(a[11]), .Y(n145) );
  AOI222XL U318 ( .A0(n148), .A1(n329), .B0(n275), .B1(n147), .C0(n146), .C1(
        n296), .Y(n151) );
  OAI21XL U319 ( .A0(n234), .A1(n190), .B0(n241), .Y(n280) );
  AOI2BB2X1 U320 ( .B0(b[2]), .B1(n158), .A0N(b[2]), .A1N(n157), .Y(n303) );
  OAI21XL U321 ( .A0(a[1]), .A1(n332), .B0(n331), .Y(n179) );
  OAI22XL U322 ( .A0(n213), .A1(n162), .B0(n214), .B1(n161), .Y(n163) );
  OAI22XL U323 ( .A0(a[1]), .A1(n170), .B0(a[2]), .B1(n215), .Y(n171) );
  OAI21XL U324 ( .A0(a[4]), .A1(n214), .B0(n172), .Y(n173) );
  OAI21XL U325 ( .A0(n252), .A1(n42), .B0(n173), .Y(n183) );
  OAI22XL U326 ( .A0(n305), .A1(n183), .B0(n253), .B1(n174), .Y(n175) );
  OAI221XL U327 ( .A0(b[1]), .A1(n332), .B0(n190), .B1(n321), .C0(n331), .Y(
        n177) );
  OAI21XL U328 ( .A0(n181), .A1(n42), .B0(n180), .Y(n347) );
  OAI21XL U329 ( .A0(b[3]), .A1(n183), .B0(n182), .Y(n184) );
  OAI21XL U330 ( .A0(n215), .A1(n282), .B0(n188), .Y(n276) );
  OAI22XL U331 ( .A0(n284), .A1(n342), .B0(n276), .B1(n283), .Y(n206) );
  AOI222XL U332 ( .A0(n251), .A1(n193), .B0(n192), .B1(n191), .C0(n190), .C1(
        n189), .Y(n197) );
  OAI22XL U333 ( .A0(n197), .A1(n195), .B0(n255), .B1(n194), .Y(n205) );
  OAI21XL U334 ( .A0(a[2]), .A1(n332), .B0(n331), .Y(n203) );
  OAI221XL U335 ( .A0(b[2]), .A1(n332), .B0(n42), .B1(n321), .C0(n331), .Y(
        n196) );
  OAI22XL U336 ( .A0(n197), .A1(n326), .B0(n324), .B1(n276), .Y(n198) );
  AO22X1 U337 ( .A0(n298), .A1(n201), .B0(n313), .B1(n200), .Y(n202) );
  OAI21XL U338 ( .A0(b[3]), .A1(n332), .B0(n331), .Y(n224) );
  OAI22XL U339 ( .A0(n213), .A1(n322), .B0(n214), .B1(n207), .Y(n208) );
  OAI22XL U340 ( .A0(a[4]), .A1(n215), .B0(a[6]), .B1(n214), .Y(n216) );
  OAI22XL U341 ( .A0(n295), .A1(n42), .B0(n217), .B1(n216), .Y(n227) );
  OAI22XL U342 ( .A0(n284), .A1(n218), .B0(n305), .B1(n227), .Y(n219) );
  AOI221XL U343 ( .A0(n272), .A1(a[3]), .B0(n41), .B1(n221), .C0(n317), .Y(
        n222) );
  OAI21XL U344 ( .A0(b[3]), .A1(n227), .B0(n226), .Y(n228) );
  OAI21XL U345 ( .A0(a[4]), .A1(n332), .B0(n331), .Y(n237) );
  OAI22XL U346 ( .A0(n300), .A1(n232), .B0(n238), .B1(n326), .Y(n233) );
  OAI221XL U347 ( .A0(b[4]), .A1(n332), .B0(n234), .B1(n321), .C0(n331), .Y(
        n235) );
  OAI2BB2XL U348 ( .B0(n42), .B1(n239), .A0N(n42), .A1N(n238), .Y(n247) );
  OAI221XL U349 ( .A0(a[5]), .A1(n332), .B0(n251), .B1(n321), .C0(n331), .Y(
        n261) );
  OAI2BB2XL U350 ( .B0(b[2]), .B1(n267), .A0N(b[2]), .A1N(n264), .Y(n258) );
  OAI22XL U351 ( .A0(n256), .A1(n255), .B0(n254), .B1(n253), .Y(n257) );
  OAI21XL U352 ( .A0(b[5]), .A1(n332), .B0(n331), .Y(n259) );
  OAI221XL U353 ( .A0(a[7]), .A1(n332), .B0(n282), .B1(n321), .C0(n331), .Y(
        n291) );
  OAI22XL U354 ( .A0(n285), .A1(n284), .B0(n294), .B1(n283), .Y(n286) );
  OAI21XL U355 ( .A0(b[7]), .A1(n332), .B0(n331), .Y(n289) );
  AOI2BB2X1 U356 ( .B0(n296), .B1(n295), .A0N(n324), .A1N(n294), .Y(n297) );
  OAI21XL U357 ( .A0(b[8]), .A1(n332), .B0(n331), .Y(n304) );
  AOI222XL U358 ( .A0(n308), .A1(n307), .B0(n308), .B1(n306), .C0(n307), .C1(
        n305), .Y(n320) );
  OAI222XL U359 ( .A0(n314), .A1(n324), .B0(n313), .B1(n312), .C0(n326), .C1(
        n311), .Y(n319) );
  OAI22XL U360 ( .A0(a[8]), .A1(n332), .B0(n315), .B1(n321), .Y(n316) );
  OAI21XL U361 ( .A0(n317), .A1(n316), .B0(b[8]), .Y(n318) );
  OAI221XL U362 ( .A0(a[9]), .A1(n332), .B0(n322), .B1(n321), .C0(n331), .Y(
        n335) );
  OAI22XL U363 ( .A0(n326), .A1(n325), .B0(n324), .B1(n323), .Y(n327) );
  AOI221XL U364 ( .A0(n330), .A1(n329), .B0(n328), .B1(n329), .C0(n327), .Y(
        n334) );
  OAI21XL U365 ( .A0(b[9]), .A1(n332), .B0(n331), .Y(n333) );
endmodule
